module NN(
    input clk,
    input a,
    output logic b
);

always_ff @( posedge clk )
begin:

end



endmodule